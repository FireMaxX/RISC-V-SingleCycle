
module instructionmemory#(
    parameter INS_ADDRESS = 9,
    parameter INS_W = 32
     )(
    input logic [ INS_ADDRESS -1:0] ra , // Read address of the instruction memory , comes from PC
    output logic [ INS_W -1:0] rd // Read Data
    );
    

logic [INS_W-1 :0] Inst_mem [(2**(INS_ADDRESS-2))-1:0];

assign Inst_mem[0 ]=32'b00000000000000000000000000010011;//			#r0 =0		(r0=0)
assign Inst_mem[1 ]=32'b00000000100000000000000010010011;//			#r1 =r0+8	(r1=8)
assign Inst_mem[2 ]=32'b00000000010000000000000100010011;//			#r2 =r0+4	(r2=4)
assign Inst_mem[3 ]=32'b00000000001000001110000110110011;//			#r3 =r1|r2	(r3=12)
assign Inst_mem[4 ]=32'b00000000000000010110001000110011;//			#r4 =r2|r0	(r4=4)

assign Inst_mem[5 ]=32'b00000000001000001000011001100011;//			#if $r1=r2 then pc=pc+12	(r1!=r2, not jump
assign Inst_mem[6 ]=32'b00000000100000000000000100010011;// 		#r2 = r2+4					(r2=8)
assign Inst_mem[7 ]=32'b00000000001000001000010001100011;// 		#if $r1=r2 then pc=pc+8		(r1=r2, jump)
assign Inst_mem[8 ]=32'b00000000000100001010000000100011;// 		#M[r1+0] = r1	(M[8]=8)	if(M[8]!=0), BEQ 
assign Inst_mem[9 ]=32'b00000000001000001010000010100011;// 		#M[r1+1] = r2	(M[9]=8)	if(M[9]=8), BEQ 

assign Inst_mem[10]=32'b00000000010000000000000100010011;// 		#r2 =r0+4	(r2=4) 

assign Inst_mem[11]=32'b00000000010000010001011001100011;// 		#if $r2!=r4 then pc=pc+12	(r2=r4, not jump)
assign Inst_mem[12]=32'b00000000100000000000000110010011;// 		#r3 =r0+8	(r3=8)
assign Inst_mem[13]=32'b00000000001000001001010001100011;// 		#if $r1!=r2 then pc=pc+8	(r1!=r2, jump)
assign Inst_mem[14]=32'b00000000001100001010000100100011;// 		#M[r1+2] = r3	(M[10]=12)	if(M[10]!=0), bne
assign Inst_mem[15]=32'b00000000001100001010000110100011;// 		#M[r1+3] = r3	(M[11]=8)	if(M[11]=8),  bne

assign Inst_mem[16]=32'b00000000010000000000000100010011;// 		#r2 =r0+4	(r2=4)
assign Inst_mem[17]=32'b00000000110000000000000110010011;// 		#r3 =r0+8	(r3=12)	

assign Inst_mem[18]=32'b00000000001000001100011001100011;// 		#if(r1<r2) then pc=pc+12	(r1>r2, not jump)
assign Inst_mem[19]=32'b00000000100000000000000110010011;// 		#r3 =r0+8	(r3=8)
assign Inst_mem[20]=32'b00000000000100010100010001100011;// 		#if(r2<r1) then pc=pc+12	(r2<r1, jump)
assign Inst_mem[21]=32'b00000000001100001010001000100011;// 		#M[r1+4] = r3	(M[12]=12)	if(M[12]!=0), blt
assign Inst_mem[22]=32'b00000000001100001010001010100011;// 		#M[r1+5] = r3	(M[13]=8)	if(M[13]=8),  blt

assign Inst_mem[23]=32'b00000000010000000000000100010011;// 		#r2 =r0+4	(r2=4)
assign Inst_mem[24]=32'b00000000110000000000000110010011;// 		#r3 =r0+8	(r3=12)	

assign Inst_mem[25]=32'b00000000000100010101011001100011;// 		#if(r2>r1) then pc=pc+12	(r1>r2, not jump)
assign Inst_mem[26]=32'b00000000100000000000000110010011;// 		#r3 =r0+8	(r3=8)
assign Inst_mem[27]=32'b00000000001000001101010001100011;// 		#if(r1>r2) then pc=pc+8	(r1>r2, jump)
assign Inst_mem[28]=32'b00000000001100001010001100100011;// 		#M[r1+6] = r3	(M[14]=12)	if(M[14]!=0), bge
assign Inst_mem[29]=32'b00000000001100001010001110100011;// 		#M[r1+7] = r3	(M[15]=8)	if(M[15]=8),  bge

assign Inst_mem[30]=32'b11111111110000000000000100010011;// 		#r2 =r0+4	(r2=-4)
assign Inst_mem[31]=32'b00000000110000000000000110010011;// 		#r3 =r0+8	(r3=12)	

assign Inst_mem[32]=32'b00000000000100010110011001100011;// 		#if(r2<r1) then pc=pc+12	(r2>r1, not jump)
assign Inst_mem[33]=32'b00000000100000000000000110010011;// 		#r3 =r0+8	(r3=8)
assign Inst_mem[34]=32'b00000000001000001110010001100011;// 		#if(r1<r2) then pc=pc+8	(r1<r2, jump)
assign Inst_mem[35]=32'b00000000001100001010010000100011;// 		#M[r1+8] = r3	(M[16]=12)	if(M[16]!=0), blt
assign Inst_mem[36]=32'b00000000001100001010010010100011;// 		#M[r1+9] = r3	(M[17]=8)	if(M[17]=8),  blt

assign Inst_mem[37]=32'b00000000110000000000000110010011;// 		#r3 =r0+8	(r3=12)	

assign Inst_mem[38]=32'b00000000001000001111011001100011;// 		#if(r1>r2) then pc=pc+12	(r1<r2, not jump)
assign Inst_mem[39]=32'b00000000100000000000000110010011;// 		#r3 =r0+8	(r3=8)
assign Inst_mem[40]=32'b00000000000100010111010001100011;// 		#if(r2>r1) then pc=pc+8		(r1<r2, jump)
assign Inst_mem[41]=32'b00000000001100001010010100100011;// 		#M[r1+10] = r3	(M[18]=12)	if(M[18]!=0), bge
assign Inst_mem[42]=32'b00000000001100001010010110100011;// 		#M[r1+11] = r3	(M[19]=8)	if(M[19]=8),  bge

assign Inst_mem[43]=32'b00000000010000000000000100010011;// 		#r2 =r0+4	(r2=4)
assign Inst_mem[44]=32'b00000000110000000000000110010011;// 		#r3 =r0+8	(r3=12)	

assign Inst_mem[45]=32'b00000000100000000000001011101111;// 		#jump to PC+8, r5=pc+4
assign Inst_mem[46]=32'b00000000100000000000000110010011;// 		#r3 =r0+8	(r3=8)
assign Inst_mem[47]=32'b00000000001100001010011000100011;// 		#M[r1+12] = r3	(M[20]=12)	if(M[20]=12),  ja

assign Inst_mem[48]=32'b00000000110000000000000110010011;// 		#r3 =r0+8	(r3=12)	

assign Inst_mem[49]=32'b00001100110000000000001101100111;// 		#jump to (51+0)^2, r6=pc+4   **
assign Inst_mem[50]=32'b00000000100000000000000110010011;// 		#r3 =r0+8	(r3=8)
assign Inst_mem[51]=32'b00000000001100001010011010100011;// 		#M[r1+13] = r3	(M[21]=12)	if(M[21]=12),  ja

assign Inst_mem[52]=32'b00000000000000000001001110110111;// 		#r7=00001000
assign Inst_mem[53]=32'b00000000011100001010011100100011;// 		#M[r1+14] = r7	(M[22]=r7)	 lu

assign Inst_mem[54]=32'b00000000000000000001010000010111;// 		#r8=54^2+00001000=000010D8
assign Inst_mem[55]=32'b00000000100000001010011110100011;// 		#M[r1+15] = r8	(M[23]=r8)	if(M[22]=r8),  auipc

assign Inst_mem[56]=32'b00000000110000000000000110010011;// 		#r3 =r0+8	(r3=12)
	//**********************
assign Inst_mem[57]=32'b00000000000000000000010100000011;// 		#R10=M[0]		r10=8
assign Inst_mem[58]=32'b00000000000100000000010110000011;// 		#R11=M[1]		r11=FFFFFFF8
assign Inst_mem[59]=32'b00000000001000000001011000000011;// 		#R12=M[2]		r12=00007FFF
assign Inst_mem[60]=32'b00000000001100000001011010000011;// 		#R13=M[3]		r13=FFFFFFFF
assign Inst_mem[61]=32'b00000000000000000100011100000011;// 		#R14=M[0]		r14=8
assign Inst_mem[62]=32'b00000000000100000100011110000011;// 		#R15=M[1]		r15=000000F8
assign Inst_mem[63]=32'b00000000001000000101100000000011;// 		#R16=M[2]		r16=00007FFF
assign Inst_mem[64]=32'b00000000001100000101100010000011;// 		#R17=M[3]		r17=0000FFFF
//*********************
assign Inst_mem[65]=32'b11111111110000000000010010010011;// 		#r9 =r0-4		(r9=-4)

assign Inst_mem[66]=32'b00000000010000000000110000100011;// 		#M[0+24]=r4		(M[0+24]=4)                                   
assign Inst_mem[67]=32'b00000000100100000000110010100011;// 		#M[0+25]=r9		(M[0+25]=FFFFFFFC)
assign Inst_mem[68]=32'b00000000010000000001110100100011;// 		#M[0+26]=r4		(M[0+26]=4)
assign Inst_mem[69]=32'b00000000100100000001110110100011;// 		#M[0+27]=r9		(M[0+27]=FFFFFFFC)

assign Inst_mem[70]=32'b00000000001000000000001000010011;// 		#r4 =r0+2		(r4=2)
assign Inst_mem[71]=32'b11111111111000000000001010010011;// 		#r5 =r0-2		(r5=-2)

assign Inst_mem[72]=32'b00000000010000001001100100110011;// 		#R18=R1<<R4 	(R18 = 8<<2)	R18=0000020
assign Inst_mem[73]=32'b00000000010000101101100110110011;// 		#R19=R5>>R4		(R19 = -2>>2) 	R19=3FFFFFF
assign Inst_mem[74]=32'b01000000010000101101101000110011;// 		#R20=R5>>>R4	(R20 = -2>>2)	R20=FFFFFFF

assign Inst_mem[75]=32'b00000000001000001010101010110011;// 		#if R1<R2, R21=1	(R21=0)
assign Inst_mem[76]=32'b00000000000100010010101100110011;// 		#if R2<R1, R22=1	(R22=1)
assign Inst_mem[77]=32'b00000000000100101011101110110011;// 		#if R5<R1, R23=1	(R23=0)
assign Inst_mem[78]=32'b00000000010100001011110000110011;// 		#if R1<R5, R24=1	(R24=1)
assign Inst_mem[79]=32'b00000000100000001010110010010011;// 		#if R1<8,  R25=1	(R25=0)
assign Inst_mem[80]=32'b00000001000000001010110100010011;// 		#if R1<16, R26=1	(R26=1)

assign Inst_mem[81]=32'b11111111110000000000001010010011;// 		#r5 =r0-4		(r5=-4)

assign Inst_mem[82]=32'b11111111111000001011110110010011;// 		#if R1<u(-2),  R27=1	(R27=1)
assign Inst_mem[83]=32'b11111111111000101011111000010011;// 		#if R5<u(-2),  R28=1	(R28=1)

assign Inst_mem[84]=32'b00000000000100101001111010010011;// 		#R29=R5<<1 	(R29=FFFFFFF8)
assign Inst_mem[85]=32'b00000000000100101101111100010011;// 		#R30=R5>>1 	(R30=7FFFFFFE)
assign Inst_mem[86]=32'b01000000000100101101111110010011;// 		#R31=R5>>1	(R31=FFFFFFFE)	**** i add inst[30]=1

assign Inst_mem[87]=32'b00000000101000001100001100010011;// 		#R6=R1 xor A	(R6=00000002)
assign Inst_mem[88]=32'b00000000001000001110001110010011;// 		#R7=R1 or 2		(R7=0000000A)
assign Inst_mem[89]=32'b00000000101000001111010000010011;// 		#R8=R1 and A	(R8=00000008)
assign Inst_mem[90]=32'b00000000001000001100010010110011;// 		#R9=R1 or R2	(R9=0000000C)


assign rd =  Inst_mem [ra[INS_ADDRESS-1:2]];  

//      genvar i;
//      generate
//          for (i = 15; i < 127; i++) begin
//              assign Inst_mem[i] = 32'h00007033;
//          end
//      endgenerate

endmodule